VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Maj_opamp
  CLASS BLOCK ;
  FOREIGN tt_um_Maj_opamp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.751700 ;
    PORT
      LAYER li1 ;
        RECT 106.400 21.020 106.570 26.060 ;
        RECT 107.980 21.020 108.150 26.060 ;
        RECT 109.560 21.020 109.730 26.060 ;
        RECT 105.440 12.210 105.610 16.160 ;
        RECT 107.020 12.210 107.190 16.160 ;
        RECT 108.600 12.210 108.770 16.160 ;
      LAYER mcon ;
        RECT 106.400 25.795 106.570 25.965 ;
        RECT 106.400 25.435 106.570 25.605 ;
        RECT 106.400 25.075 106.570 25.245 ;
        RECT 106.400 24.715 106.570 24.885 ;
        RECT 106.400 24.355 106.570 24.525 ;
        RECT 106.400 23.995 106.570 24.165 ;
        RECT 106.400 23.635 106.570 23.805 ;
        RECT 106.400 23.275 106.570 23.445 ;
        RECT 106.400 22.915 106.570 23.085 ;
        RECT 106.400 22.555 106.570 22.725 ;
        RECT 106.400 22.195 106.570 22.365 ;
        RECT 106.400 21.835 106.570 22.005 ;
        RECT 106.400 21.475 106.570 21.645 ;
        RECT 106.400 21.115 106.570 21.285 ;
        RECT 107.980 25.795 108.150 25.965 ;
        RECT 107.980 25.435 108.150 25.605 ;
        RECT 107.980 25.075 108.150 25.245 ;
        RECT 107.980 24.715 108.150 24.885 ;
        RECT 107.980 24.355 108.150 24.525 ;
        RECT 107.980 23.995 108.150 24.165 ;
        RECT 107.980 23.635 108.150 23.805 ;
        RECT 107.980 23.275 108.150 23.445 ;
        RECT 107.980 22.915 108.150 23.085 ;
        RECT 107.980 22.555 108.150 22.725 ;
        RECT 107.980 22.195 108.150 22.365 ;
        RECT 107.980 21.835 108.150 22.005 ;
        RECT 107.980 21.475 108.150 21.645 ;
        RECT 107.980 21.115 108.150 21.285 ;
        RECT 109.560 25.795 109.730 25.965 ;
        RECT 109.560 25.435 109.730 25.605 ;
        RECT 109.560 25.075 109.730 25.245 ;
        RECT 109.560 24.715 109.730 24.885 ;
        RECT 109.560 24.355 109.730 24.525 ;
        RECT 109.560 23.995 109.730 24.165 ;
        RECT 109.560 23.635 109.730 23.805 ;
        RECT 109.560 23.275 109.730 23.445 ;
        RECT 109.560 22.915 109.730 23.085 ;
        RECT 109.560 22.555 109.730 22.725 ;
        RECT 109.560 22.195 109.730 22.365 ;
        RECT 109.560 21.835 109.730 22.005 ;
        RECT 109.560 21.475 109.730 21.645 ;
        RECT 109.560 21.115 109.730 21.285 ;
        RECT 105.440 15.900 105.610 16.070 ;
        RECT 105.440 15.540 105.610 15.710 ;
        RECT 105.440 15.180 105.610 15.350 ;
        RECT 105.440 14.820 105.610 14.990 ;
        RECT 105.440 14.460 105.610 14.630 ;
        RECT 105.440 14.100 105.610 14.270 ;
        RECT 105.440 13.740 105.610 13.910 ;
        RECT 105.440 13.380 105.610 13.550 ;
        RECT 105.440 13.020 105.610 13.190 ;
        RECT 105.440 12.660 105.610 12.830 ;
        RECT 105.440 12.300 105.610 12.470 ;
        RECT 107.020 15.900 107.190 16.070 ;
        RECT 107.020 15.540 107.190 15.710 ;
        RECT 107.020 15.180 107.190 15.350 ;
        RECT 107.020 14.820 107.190 14.990 ;
        RECT 107.020 14.460 107.190 14.630 ;
        RECT 107.020 14.100 107.190 14.270 ;
        RECT 107.020 13.740 107.190 13.910 ;
        RECT 107.020 13.380 107.190 13.550 ;
        RECT 107.020 13.020 107.190 13.190 ;
        RECT 107.020 12.660 107.190 12.830 ;
        RECT 107.020 12.300 107.190 12.470 ;
        RECT 108.600 15.900 108.770 16.070 ;
        RECT 108.600 15.540 108.770 15.710 ;
        RECT 108.600 15.180 108.770 15.350 ;
        RECT 108.600 14.820 108.770 14.990 ;
        RECT 108.600 14.460 108.770 14.630 ;
        RECT 108.600 14.100 108.770 14.270 ;
        RECT 108.600 13.740 108.770 13.910 ;
        RECT 108.600 13.380 108.770 13.550 ;
        RECT 108.600 13.020 108.770 13.190 ;
        RECT 108.600 12.660 108.770 12.830 ;
        RECT 108.600 12.300 108.770 12.470 ;
      LAYER met1 ;
        RECT 106.370 24.910 106.600 26.040 ;
        RECT 107.950 24.910 108.180 26.040 ;
        RECT 109.530 24.910 109.760 26.040 ;
        RECT 106.370 24.760 106.700 24.910 ;
        RECT 106.370 22.750 106.810 24.760 ;
        RECT 106.370 21.040 106.600 22.750 ;
        RECT 107.950 22.690 108.270 24.910 ;
        RECT 109.530 22.690 109.850 24.910 ;
        RECT 107.950 21.040 108.180 22.690 ;
        RECT 109.530 21.040 109.760 22.690 ;
        RECT 105.410 15.520 105.640 16.140 ;
        RECT 106.990 15.540 107.220 16.140 ;
        RECT 108.570 15.550 108.800 16.140 ;
        RECT 105.410 13.300 105.810 15.520 ;
        RECT 106.990 13.320 107.400 15.540 ;
        RECT 108.570 13.330 108.980 15.550 ;
        RECT 105.410 12.230 105.640 13.300 ;
        RECT 106.990 12.230 107.220 13.320 ;
        RECT 108.570 12.230 108.800 13.330 ;
      LAYER via ;
        RECT 106.405 24.540 106.665 24.800 ;
        RECT 106.405 24.220 106.665 24.480 ;
        RECT 106.405 23.900 106.665 24.160 ;
        RECT 106.405 23.580 106.665 23.840 ;
        RECT 106.405 23.260 106.665 23.520 ;
        RECT 106.405 22.940 106.665 23.200 ;
        RECT 107.990 24.445 108.250 24.705 ;
        RECT 107.990 24.125 108.250 24.385 ;
        RECT 107.990 23.805 108.250 24.065 ;
        RECT 107.990 23.485 108.250 23.745 ;
        RECT 107.990 23.165 108.250 23.425 ;
        RECT 107.990 22.845 108.250 23.105 ;
        RECT 109.570 24.435 109.830 24.695 ;
        RECT 109.570 24.115 109.830 24.375 ;
        RECT 109.570 23.795 109.830 24.055 ;
        RECT 109.570 23.475 109.830 23.735 ;
        RECT 109.570 23.155 109.830 23.415 ;
        RECT 109.570 22.835 109.830 23.095 ;
        RECT 105.435 15.155 105.695 15.415 ;
        RECT 105.435 14.835 105.695 15.095 ;
        RECT 105.435 14.515 105.695 14.775 ;
        RECT 105.435 14.195 105.695 14.455 ;
        RECT 105.435 13.875 105.695 14.135 ;
        RECT 105.435 13.555 105.695 13.815 ;
        RECT 107.015 15.145 107.275 15.405 ;
        RECT 107.015 14.825 107.275 15.085 ;
        RECT 107.015 14.505 107.275 14.765 ;
        RECT 107.015 14.185 107.275 14.445 ;
        RECT 107.015 13.865 107.275 14.125 ;
        RECT 107.015 13.545 107.275 13.805 ;
        RECT 108.605 15.135 108.865 15.395 ;
        RECT 108.605 14.815 108.865 15.075 ;
        RECT 108.605 14.495 108.865 14.755 ;
        RECT 108.605 14.175 108.865 14.435 ;
        RECT 108.605 13.855 108.865 14.115 ;
        RECT 108.605 13.535 108.865 13.795 ;
      LAYER met2 ;
        RECT 106.120 22.990 109.910 24.910 ;
        RECT 106.120 22.690 114.850 22.990 ;
        RECT 106.750 21.390 114.850 22.690 ;
        RECT 106.780 15.630 108.430 21.390 ;
        RECT 105.070 13.160 109.210 15.630 ;
      LAYER via2 ;
        RECT 112.660 21.650 114.540 22.730 ;
      LAYER met3 ;
        RECT 112.300 21.390 114.850 22.990 ;
      LAYER via3 ;
        RECT 112.640 21.630 114.560 22.750 ;
      LAYER met4 ;
        RECT 118.245 22.990 147.855 43.895 ;
        RECT 112.300 21.390 147.855 22.990 ;
        RECT 113.170 8.590 114.070 21.390 ;
        RECT 118.245 14.285 147.855 21.390 ;
        RECT 113.170 7.690 152.710 8.590 ;
        RECT 151.810 0.000 152.710 7.690 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.500000 ;
    PORT
      LAYER li1 ;
        RECT 101.790 21.560 102.290 21.730 ;
        RECT 101.790 18.010 102.290 18.180 ;
      LAYER mcon ;
        RECT 101.955 21.560 102.125 21.730 ;
        RECT 101.955 18.010 102.125 18.180 ;
      LAYER met1 ;
        RECT 101.520 21.520 102.530 21.980 ;
        RECT 101.810 17.980 102.270 18.210 ;
      LAYER via ;
        RECT 101.570 21.520 102.480 21.980 ;
      LAYER met2 ;
        RECT 101.570 21.470 102.480 22.030 ;
      LAYER via2 ;
        RECT 101.570 21.520 102.480 21.980 ;
      LAYER met3 ;
        RECT 101.520 21.495 102.530 22.005 ;
      LAYER via3 ;
        RECT 101.570 21.520 102.480 21.980 ;
      LAYER met4 ;
        RECT 101.565 21.515 102.485 21.985 ;
        RECT 101.570 4.230 102.470 21.515 ;
        RECT 101.570 3.200 133.390 4.230 ;
        RECT 132.490 0.000 133.390 3.200 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.500000 ;
    PORT
      LAYER li1 ;
        RECT 99.335 21.560 99.835 21.730 ;
        RECT 99.335 18.010 99.835 18.180 ;
      LAYER mcon ;
        RECT 99.500 21.560 99.670 21.730 ;
        RECT 99.500 18.010 99.670 18.180 ;
      LAYER met1 ;
        RECT 99.040 21.520 100.030 21.940 ;
        RECT 99.355 17.980 99.815 18.210 ;
      LAYER via ;
        RECT 99.090 21.520 99.980 21.940 ;
      LAYER met2 ;
        RECT 99.090 21.470 99.980 21.990 ;
      LAYER via2 ;
        RECT 99.090 21.520 99.980 21.940 ;
      LAYER met3 ;
        RECT 99.040 21.495 100.030 21.965 ;
      LAYER via3 ;
        RECT 99.090 21.520 99.980 21.940 ;
      LAYER met4 ;
        RECT 99.080 21.945 99.980 22.090 ;
        RECT 99.080 21.515 99.985 21.945 ;
        RECT 99.080 2.340 99.980 21.515 ;
        RECT 99.080 1.440 114.070 2.340 ;
        RECT 113.170 0.000 114.070 1.440 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.610 0.100 94.750 1.000 ;
        RECT 93.850 0.000 94.750 0.100 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.250 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.250 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 100.800 26.765 103.260 26.780 ;
        RECT 98.385 22.590 103.260 26.765 ;
        RECT 98.385 22.575 100.845 22.590 ;
        RECT 104.860 19.940 110.480 26.780 ;
      LAYER li1 ;
        RECT 96.120 28.290 96.810 30.450 ;
        RECT 97.900 27.240 115.800 28.590 ;
        RECT 99.350 26.585 99.850 27.240 ;
        RECT 100.450 26.600 101.150 26.640 ;
        RECT 101.800 26.600 102.300 27.240 ;
        RECT 107.600 26.600 108.100 27.240 ;
        RECT 100.450 26.590 103.080 26.600 ;
        RECT 100.400 26.585 103.080 26.590 ;
        RECT 98.565 26.440 103.080 26.585 ;
        RECT 98.565 26.415 100.665 26.440 ;
        RECT 98.565 25.690 98.735 26.415 ;
        RECT 98.550 25.340 99.350 25.690 ;
        RECT 98.565 22.925 98.735 25.340 ;
        RECT 99.135 23.650 99.305 25.340 ;
        RECT 100.495 22.925 100.665 26.415 ;
        RECT 98.565 22.755 100.665 22.925 ;
        RECT 100.980 26.430 103.080 26.440 ;
        RECT 100.980 22.940 101.150 26.430 ;
        RECT 102.340 25.690 102.510 25.705 ;
        RECT 102.910 25.690 103.080 26.430 ;
        RECT 105.040 26.430 110.300 26.600 ;
        RECT 105.040 25.690 105.210 26.430 ;
        RECT 105.580 25.710 105.810 26.430 ;
        RECT 107.160 25.710 107.390 26.430 ;
        RECT 108.740 25.710 108.970 26.430 ;
        RECT 102.290 25.240 105.210 25.690 ;
        RECT 102.340 23.665 102.510 25.240 ;
        RECT 102.910 22.940 103.080 25.240 ;
        RECT 100.980 22.770 103.080 22.940 ;
        RECT 105.040 20.290 105.210 25.240 ;
        RECT 105.610 21.020 105.780 25.710 ;
        RECT 107.190 21.020 107.360 25.710 ;
        RECT 108.770 21.020 108.940 25.710 ;
        RECT 110.130 20.290 110.300 26.430 ;
        RECT 105.040 20.120 110.300 20.290 ;
      LAYER mcon ;
        RECT 96.200 28.380 96.730 30.350 ;
        RECT 98.725 28.315 98.895 28.485 ;
        RECT 103.730 27.635 104.260 28.165 ;
        RECT 99.135 25.305 99.305 25.475 ;
        RECT 99.135 24.945 99.305 25.115 ;
        RECT 99.135 24.585 99.305 24.755 ;
        RECT 99.135 24.225 99.305 24.395 ;
        RECT 99.135 23.865 99.305 24.035 ;
        RECT 105.610 25.795 105.780 25.965 ;
        RECT 107.190 25.795 107.360 25.965 ;
        RECT 108.770 25.795 108.940 25.965 ;
        RECT 102.340 25.320 102.510 25.490 ;
        RECT 102.340 24.960 102.510 25.130 ;
        RECT 102.340 24.600 102.510 24.770 ;
        RECT 102.340 24.240 102.510 24.410 ;
        RECT 102.340 23.880 102.510 24.050 ;
        RECT 105.610 25.435 105.780 25.605 ;
        RECT 105.610 25.075 105.780 25.245 ;
        RECT 105.610 24.715 105.780 24.885 ;
        RECT 105.610 24.355 105.780 24.525 ;
        RECT 105.610 23.995 105.780 24.165 ;
        RECT 105.610 23.635 105.780 23.805 ;
        RECT 105.610 23.275 105.780 23.445 ;
        RECT 105.610 22.915 105.780 23.085 ;
        RECT 105.610 22.555 105.780 22.725 ;
        RECT 105.610 22.195 105.780 22.365 ;
        RECT 105.610 21.835 105.780 22.005 ;
        RECT 105.610 21.475 105.780 21.645 ;
        RECT 105.610 21.115 105.780 21.285 ;
        RECT 107.190 25.435 107.360 25.605 ;
        RECT 107.190 25.075 107.360 25.245 ;
        RECT 107.190 24.715 107.360 24.885 ;
        RECT 107.190 24.355 107.360 24.525 ;
        RECT 107.190 23.995 107.360 24.165 ;
        RECT 107.190 23.635 107.360 23.805 ;
        RECT 107.190 23.275 107.360 23.445 ;
        RECT 107.190 22.915 107.360 23.085 ;
        RECT 107.190 22.555 107.360 22.725 ;
        RECT 107.190 22.195 107.360 22.365 ;
        RECT 107.190 21.835 107.360 22.005 ;
        RECT 107.190 21.475 107.360 21.645 ;
        RECT 107.190 21.115 107.360 21.285 ;
        RECT 108.770 25.435 108.940 25.605 ;
        RECT 108.770 25.075 108.940 25.245 ;
        RECT 108.770 24.715 108.940 24.885 ;
        RECT 108.770 24.355 108.940 24.525 ;
        RECT 108.770 23.995 108.940 24.165 ;
        RECT 108.770 23.635 108.940 23.805 ;
        RECT 108.770 23.275 108.940 23.445 ;
        RECT 108.770 22.915 108.940 23.085 ;
        RECT 108.770 22.555 108.940 22.725 ;
        RECT 108.770 22.195 108.940 22.365 ;
        RECT 108.770 21.835 108.940 22.005 ;
        RECT 108.770 21.475 108.940 21.645 ;
        RECT 108.770 21.115 108.940 21.285 ;
      LAYER met1 ;
        RECT 1.220 43.960 2.820 46.310 ;
        RECT 1.220 42.380 104.820 43.960 ;
        RECT 1.220 42.370 101.890 42.380 ;
        RECT 1.220 38.400 2.820 42.370 ;
        RECT 96.170 28.590 96.760 30.420 ;
        RECT 96.100 28.270 99.950 28.590 ;
        RECT 97.750 28.260 99.950 28.270 ;
        RECT 103.240 27.240 104.820 42.380 ;
        RECT 99.105 23.670 99.335 25.670 ;
        RECT 102.310 23.685 102.540 25.685 ;
        RECT 105.580 21.040 105.810 26.040 ;
        RECT 107.160 21.040 107.390 26.040 ;
        RECT 108.740 21.040 108.970 26.040 ;
      LAYER via ;
        RECT 1.250 38.430 2.790 46.280 ;
      LAYER met2 ;
        RECT 1.170 38.350 2.870 46.360 ;
      LAYER via2 ;
        RECT 1.220 38.400 2.820 46.310 ;
      LAYER met3 ;
        RECT 1.170 38.350 2.870 46.370 ;
      LAYER via3 ;
        RECT 1.200 38.380 2.840 46.340 ;
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 95.340 30.800 97.590 31.230 ;
        RECT 95.340 7.240 95.770 30.800 ;
        RECT 97.160 7.240 97.590 30.800 ;
        RECT 98.405 17.370 100.765 22.370 ;
        RECT 100.860 17.370 103.220 22.370 ;
        RECT 104.450 19.200 117.310 19.630 ;
        RECT 104.450 18.170 104.880 19.200 ;
        RECT 116.880 18.170 117.310 19.200 ;
        RECT 104.450 17.740 117.310 18.170 ;
        RECT 98.450 9.090 100.810 16.780 ;
        RECT 100.900 9.090 103.260 16.780 ;
        RECT 103.950 11.540 110.260 17.140 ;
        RECT 95.340 6.810 97.590 7.240 ;
      LAYER li1 ;
        RECT 95.470 30.930 97.460 31.100 ;
        RECT 95.470 7.110 95.640 30.930 ;
        RECT 97.290 8.110 97.460 30.930 ;
        RECT 100.395 22.240 101.220 22.245 ;
        RECT 98.535 22.070 103.090 22.240 ;
        RECT 98.535 17.670 98.705 22.070 ;
        RECT 100.465 17.670 100.635 22.070 ;
        RECT 100.990 17.670 101.160 22.070 ;
        RECT 102.920 17.670 103.090 22.070 ;
        RECT 104.580 19.330 117.180 19.500 ;
        RECT 104.580 18.040 104.750 19.330 ;
        RECT 117.010 18.040 117.180 19.330 ;
        RECT 104.580 17.870 117.180 18.040 ;
        RECT 98.535 17.500 103.090 17.670 ;
        RECT 100.150 17.495 101.215 17.500 ;
        RECT 100.150 16.650 100.550 17.495 ;
        RECT 100.750 17.440 100.960 17.495 ;
        RECT 105.250 17.010 105.550 17.870 ;
        RECT 104.080 16.840 110.130 17.010 ;
        RECT 98.580 16.480 100.680 16.650 ;
        RECT 98.580 10.890 98.750 16.480 ;
        RECT 99.150 10.890 99.320 16.110 ;
        RECT 98.580 10.390 99.320 10.890 ;
        RECT 98.580 9.390 98.750 10.390 ;
        RECT 99.150 10.070 99.320 10.390 ;
        RECT 100.510 9.390 100.680 16.480 ;
        RECT 101.030 16.480 103.130 16.650 ;
        RECT 101.030 9.390 101.200 16.480 ;
        RECT 102.390 10.940 102.560 16.110 ;
        RECT 102.960 10.940 103.130 16.480 ;
        RECT 104.080 13.940 104.250 16.840 ;
        RECT 103.650 13.690 104.250 13.940 ;
        RECT 102.390 10.790 103.200 10.940 ;
        RECT 103.650 10.790 103.850 13.690 ;
        RECT 104.080 11.840 104.250 13.690 ;
        RECT 104.650 11.840 104.820 16.160 ;
        RECT 106.230 11.840 106.400 16.160 ;
        RECT 107.810 11.840 107.980 16.160 ;
        RECT 109.390 11.840 109.560 16.160 ;
        RECT 109.960 11.840 110.130 16.840 ;
        RECT 104.080 11.670 110.130 11.840 ;
        RECT 102.390 10.590 103.850 10.790 ;
        RECT 102.390 10.440 103.200 10.590 ;
        RECT 102.390 10.070 102.560 10.440 ;
        RECT 102.960 9.390 103.130 10.440 ;
        RECT 98.580 9.220 103.130 9.390 ;
        RECT 100.300 9.190 101.450 9.220 ;
        RECT 100.400 8.890 101.350 9.190 ;
        RECT 106.600 8.890 107.400 11.670 ;
        RECT 97.290 8.100 97.830 8.110 ;
        RECT 98.400 8.100 111.900 8.890 ;
        RECT 97.290 7.740 111.900 8.100 ;
        RECT 97.290 7.110 97.460 7.740 ;
        RECT 98.400 7.290 111.900 7.740 ;
        RECT 95.470 6.940 97.460 7.110 ;
      LAYER mcon ;
        RECT 99.150 15.705 99.320 15.875 ;
        RECT 99.150 15.345 99.320 15.515 ;
        RECT 99.150 14.985 99.320 15.155 ;
        RECT 99.150 14.625 99.320 14.795 ;
        RECT 99.150 14.265 99.320 14.435 ;
        RECT 99.150 13.905 99.320 14.075 ;
        RECT 99.150 13.545 99.320 13.715 ;
        RECT 99.150 13.185 99.320 13.355 ;
        RECT 99.150 12.825 99.320 12.995 ;
        RECT 99.150 12.465 99.320 12.635 ;
        RECT 99.150 12.105 99.320 12.275 ;
        RECT 99.150 11.745 99.320 11.915 ;
        RECT 99.150 11.385 99.320 11.555 ;
        RECT 99.150 11.025 99.320 11.195 ;
        RECT 99.150 10.665 99.320 10.835 ;
        RECT 99.150 10.305 99.320 10.475 ;
        RECT 102.390 15.705 102.560 15.875 ;
        RECT 102.390 15.345 102.560 15.515 ;
        RECT 102.390 14.985 102.560 15.155 ;
        RECT 102.390 14.625 102.560 14.795 ;
        RECT 102.390 14.265 102.560 14.435 ;
        RECT 102.390 13.905 102.560 14.075 ;
        RECT 102.390 13.545 102.560 13.715 ;
        RECT 102.390 13.185 102.560 13.355 ;
        RECT 102.390 12.825 102.560 12.995 ;
        RECT 102.390 12.465 102.560 12.635 ;
        RECT 102.390 12.105 102.560 12.275 ;
        RECT 102.390 11.745 102.560 11.915 ;
        RECT 102.390 11.385 102.560 11.555 ;
        RECT 102.390 11.025 102.560 11.195 ;
        RECT 102.390 10.665 102.560 10.835 ;
        RECT 104.650 15.900 104.820 16.070 ;
        RECT 104.650 15.540 104.820 15.710 ;
        RECT 104.650 15.180 104.820 15.350 ;
        RECT 104.650 14.820 104.820 14.990 ;
        RECT 104.650 14.460 104.820 14.630 ;
        RECT 104.650 14.100 104.820 14.270 ;
        RECT 104.650 13.740 104.820 13.910 ;
        RECT 104.650 13.380 104.820 13.550 ;
        RECT 104.650 13.020 104.820 13.190 ;
        RECT 104.650 12.660 104.820 12.830 ;
        RECT 104.650 12.300 104.820 12.470 ;
        RECT 106.230 15.900 106.400 16.070 ;
        RECT 106.230 15.540 106.400 15.710 ;
        RECT 106.230 15.180 106.400 15.350 ;
        RECT 106.230 14.820 106.400 14.990 ;
        RECT 106.230 14.460 106.400 14.630 ;
        RECT 106.230 14.100 106.400 14.270 ;
        RECT 106.230 13.740 106.400 13.910 ;
        RECT 106.230 13.380 106.400 13.550 ;
        RECT 106.230 13.020 106.400 13.190 ;
        RECT 106.230 12.660 106.400 12.830 ;
        RECT 106.230 12.300 106.400 12.470 ;
        RECT 107.810 15.900 107.980 16.070 ;
        RECT 107.810 15.540 107.980 15.710 ;
        RECT 107.810 15.180 107.980 15.350 ;
        RECT 107.810 14.820 107.980 14.990 ;
        RECT 107.810 14.460 107.980 14.630 ;
        RECT 107.810 14.100 107.980 14.270 ;
        RECT 107.810 13.740 107.980 13.910 ;
        RECT 107.810 13.380 107.980 13.550 ;
        RECT 107.810 13.020 107.980 13.190 ;
        RECT 107.810 12.660 107.980 12.830 ;
        RECT 107.810 12.300 107.980 12.470 ;
        RECT 109.390 15.900 109.560 16.070 ;
        RECT 109.390 15.540 109.560 15.710 ;
        RECT 109.390 15.180 109.560 15.350 ;
        RECT 109.390 14.820 109.560 14.990 ;
        RECT 109.390 14.460 109.560 14.630 ;
        RECT 109.390 14.100 109.560 14.270 ;
        RECT 109.390 13.740 109.560 13.910 ;
        RECT 109.390 13.380 109.560 13.550 ;
        RECT 109.390 13.020 109.560 13.190 ;
        RECT 109.390 12.660 109.560 12.830 ;
        RECT 109.390 12.300 109.560 12.470 ;
        RECT 102.390 10.305 102.560 10.475 ;
        RECT 98.420 7.300 111.860 8.870 ;
      LAYER met1 ;
        RECT 3.980 6.600 5.980 11.270 ;
        RECT 99.120 10.090 99.350 16.090 ;
        RECT 102.360 10.090 102.590 16.090 ;
        RECT 104.620 12.230 104.850 16.140 ;
        RECT 106.200 12.230 106.430 16.140 ;
        RECT 107.780 12.230 108.010 16.140 ;
        RECT 109.360 12.230 109.590 16.140 ;
        RECT 98.360 7.270 111.920 8.900 ;
        RECT 99.820 6.600 101.340 7.270 ;
        RECT 3.980 6.090 101.340 6.600 ;
        RECT 4.000 5.080 101.340 6.090 ;
        RECT 4.000 5.040 5.990 5.080 ;
      LAYER via ;
        RECT 4.030 6.700 5.930 11.270 ;
        RECT 4.030 6.090 5.940 6.700 ;
        RECT 4.050 5.040 5.940 6.090 ;
      LAYER met2 ;
        RECT 4.030 6.750 5.930 11.320 ;
        RECT 4.030 6.040 5.940 6.750 ;
        RECT 4.050 4.990 5.940 6.040 ;
      LAYER via2 ;
        RECT 4.030 6.700 5.930 11.270 ;
        RECT 4.030 6.090 5.940 6.700 ;
        RECT 4.050 5.040 5.940 6.090 ;
      LAYER met3 ;
        RECT 3.980 6.725 5.980 11.295 ;
        RECT 3.980 6.065 5.990 6.725 ;
        RECT 4.000 5.015 5.990 6.065 ;
      LAYER via3 ;
        RECT 4.030 6.700 5.930 11.270 ;
        RECT 4.030 6.090 5.940 6.700 ;
        RECT 4.050 5.040 5.940 6.090 ;
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 99.365 25.905 99.865 26.075 ;
        RECT 101.780 25.920 102.280 26.090 ;
        RECT 99.925 23.650 100.095 25.690 ;
        RECT 101.550 23.665 101.720 25.705 ;
        RECT 99.365 23.265 99.865 23.435 ;
        RECT 101.780 23.280 102.280 23.450 ;
        RECT 99.105 18.350 99.275 21.390 ;
        RECT 99.895 18.350 100.065 21.390 ;
        RECT 101.560 18.350 101.730 21.390 ;
        RECT 102.350 18.350 102.520 21.390 ;
        RECT 105.840 20.635 106.340 20.805 ;
        RECT 106.630 20.635 107.130 20.805 ;
        RECT 107.420 20.635 107.920 20.805 ;
        RECT 108.210 20.635 108.710 20.805 ;
        RECT 109.000 20.635 109.500 20.805 ;
        RECT 105.310 18.770 105.480 18.850 ;
        RECT 116.280 18.770 116.450 18.850 ;
        RECT 105.310 18.600 107.295 18.770 ;
        RECT 114.465 18.600 116.450 18.770 ;
        RECT 105.310 18.520 105.480 18.600 ;
        RECT 116.280 18.520 116.450 18.600 ;
        RECT 104.880 16.330 105.380 16.500 ;
        RECT 105.670 16.330 106.170 16.500 ;
        RECT 106.460 16.330 106.960 16.500 ;
        RECT 107.250 16.330 107.750 16.500 ;
        RECT 108.040 16.330 108.540 16.500 ;
        RECT 108.830 16.330 109.330 16.500 ;
        RECT 99.940 10.070 100.110 16.110 ;
        RECT 101.600 10.070 101.770 16.110 ;
        RECT 96.120 7.590 96.810 9.750 ;
        RECT 99.380 9.730 99.880 9.900 ;
        RECT 101.830 9.730 102.330 9.900 ;
      LAYER mcon ;
        RECT 99.530 25.905 99.700 26.075 ;
        RECT 101.945 25.920 102.115 26.090 ;
        RECT 99.925 25.305 100.095 25.475 ;
        RECT 99.925 24.945 100.095 25.115 ;
        RECT 99.925 24.585 100.095 24.755 ;
        RECT 99.925 24.225 100.095 24.395 ;
        RECT 99.925 23.865 100.095 24.035 ;
        RECT 101.550 25.320 101.720 25.490 ;
        RECT 101.550 24.960 101.720 25.130 ;
        RECT 101.550 24.600 101.720 24.770 ;
        RECT 101.550 24.240 101.720 24.410 ;
        RECT 101.550 23.880 101.720 24.050 ;
        RECT 99.530 23.265 99.700 23.435 ;
        RECT 101.945 23.280 102.115 23.450 ;
        RECT 99.105 21.045 99.275 21.215 ;
        RECT 99.105 20.685 99.275 20.855 ;
        RECT 99.105 20.325 99.275 20.495 ;
        RECT 99.105 19.965 99.275 20.135 ;
        RECT 99.105 19.605 99.275 19.775 ;
        RECT 99.105 19.245 99.275 19.415 ;
        RECT 99.105 18.885 99.275 19.055 ;
        RECT 99.105 18.525 99.275 18.695 ;
        RECT 99.895 21.045 100.065 21.215 ;
        RECT 99.895 20.685 100.065 20.855 ;
        RECT 99.895 20.325 100.065 20.495 ;
        RECT 99.895 19.965 100.065 20.135 ;
        RECT 99.895 19.605 100.065 19.775 ;
        RECT 99.895 19.245 100.065 19.415 ;
        RECT 99.895 18.885 100.065 19.055 ;
        RECT 99.895 18.525 100.065 18.695 ;
        RECT 101.560 21.045 101.730 21.215 ;
        RECT 101.560 20.685 101.730 20.855 ;
        RECT 101.560 20.325 101.730 20.495 ;
        RECT 101.560 19.965 101.730 20.135 ;
        RECT 101.560 19.605 101.730 19.775 ;
        RECT 101.560 19.245 101.730 19.415 ;
        RECT 101.560 18.885 101.730 19.055 ;
        RECT 101.560 18.525 101.730 18.695 ;
        RECT 102.350 21.045 102.520 21.215 ;
        RECT 102.350 20.685 102.520 20.855 ;
        RECT 106.005 20.635 106.175 20.805 ;
        RECT 106.795 20.635 106.965 20.805 ;
        RECT 107.585 20.635 107.755 20.805 ;
        RECT 108.375 20.635 108.545 20.805 ;
        RECT 109.165 20.635 109.335 20.805 ;
        RECT 102.350 20.325 102.520 20.495 ;
        RECT 102.350 19.965 102.520 20.135 ;
        RECT 102.350 19.605 102.520 19.775 ;
        RECT 102.350 19.245 102.520 19.415 ;
        RECT 102.350 18.885 102.520 19.055 ;
        RECT 102.350 18.525 102.520 18.695 ;
        RECT 105.315 18.600 105.485 18.770 ;
        RECT 105.675 18.600 105.845 18.770 ;
        RECT 106.035 18.600 106.205 18.770 ;
        RECT 106.395 18.600 106.565 18.770 ;
        RECT 106.755 18.600 106.925 18.770 ;
        RECT 107.115 18.600 107.285 18.770 ;
        RECT 114.470 18.600 114.640 18.770 ;
        RECT 114.830 18.600 115.000 18.770 ;
        RECT 115.190 18.600 115.360 18.770 ;
        RECT 115.550 18.600 115.720 18.770 ;
        RECT 115.910 18.600 116.080 18.770 ;
        RECT 116.270 18.600 116.440 18.770 ;
        RECT 105.045 16.330 105.215 16.500 ;
        RECT 105.835 16.330 106.005 16.500 ;
        RECT 106.625 16.330 106.795 16.500 ;
        RECT 107.415 16.330 107.585 16.500 ;
        RECT 108.205 16.330 108.375 16.500 ;
        RECT 108.995 16.330 109.165 16.500 ;
        RECT 99.940 15.705 100.110 15.875 ;
        RECT 99.940 15.345 100.110 15.515 ;
        RECT 99.940 14.985 100.110 15.155 ;
        RECT 99.940 14.625 100.110 14.795 ;
        RECT 99.940 14.265 100.110 14.435 ;
        RECT 99.940 13.905 100.110 14.075 ;
        RECT 99.940 13.545 100.110 13.715 ;
        RECT 99.940 13.185 100.110 13.355 ;
        RECT 99.940 12.825 100.110 12.995 ;
        RECT 99.940 12.465 100.110 12.635 ;
        RECT 99.940 12.105 100.110 12.275 ;
        RECT 99.940 11.745 100.110 11.915 ;
        RECT 99.940 11.385 100.110 11.555 ;
        RECT 99.940 11.025 100.110 11.195 ;
        RECT 99.940 10.665 100.110 10.835 ;
        RECT 99.940 10.305 100.110 10.475 ;
        RECT 101.600 15.705 101.770 15.875 ;
        RECT 101.600 15.345 101.770 15.515 ;
        RECT 101.600 14.985 101.770 15.155 ;
        RECT 101.600 14.625 101.770 14.795 ;
        RECT 101.600 14.265 101.770 14.435 ;
        RECT 101.600 13.905 101.770 14.075 ;
        RECT 101.600 13.545 101.770 13.715 ;
        RECT 101.600 13.185 101.770 13.355 ;
        RECT 101.600 12.825 101.770 12.995 ;
        RECT 101.600 12.465 101.770 12.635 ;
        RECT 101.600 12.105 101.770 12.275 ;
        RECT 101.600 11.745 101.770 11.915 ;
        RECT 101.600 11.385 101.770 11.555 ;
        RECT 101.600 11.025 101.770 11.195 ;
        RECT 101.600 10.665 101.770 10.835 ;
        RECT 101.600 10.305 101.770 10.475 ;
        RECT 99.545 9.730 99.715 9.900 ;
        RECT 101.995 9.730 102.165 9.900 ;
        RECT 96.200 7.685 96.730 9.655 ;
      LAYER met1 ;
        RECT 99.385 26.090 99.845 26.105 ;
        RECT 101.800 26.090 102.260 26.120 ;
        RECT 99.350 25.890 102.300 26.090 ;
        RECT 99.385 25.875 100.140 25.890 ;
        RECT 99.900 25.670 100.140 25.875 ;
        RECT 99.895 25.490 100.140 25.670 ;
        RECT 99.895 24.020 100.125 25.490 ;
        RECT 101.520 24.020 101.750 25.685 ;
        RECT 99.895 23.840 100.670 24.020 ;
        RECT 99.895 23.670 100.125 23.840 ;
        RECT 99.385 23.235 99.845 23.465 ;
        RECT 99.075 18.670 99.305 21.370 ;
        RECT 98.480 18.430 99.305 18.670 ;
        RECT 98.480 17.670 98.720 18.430 ;
        RECT 99.075 18.370 99.305 18.430 ;
        RECT 99.865 21.320 100.095 21.370 ;
        RECT 100.460 21.320 100.670 23.840 ;
        RECT 99.865 21.140 100.670 21.320 ;
        RECT 100.980 23.840 101.750 24.020 ;
        RECT 100.980 22.590 101.190 23.840 ;
        RECT 101.520 23.685 101.750 23.840 ;
        RECT 101.800 23.250 102.260 23.480 ;
        RECT 100.980 22.420 104.160 22.590 ;
        RECT 100.980 21.330 101.190 22.420 ;
        RECT 101.530 21.330 101.760 21.370 ;
        RECT 100.980 21.150 101.760 21.330 ;
        RECT 99.865 18.370 100.095 21.140 ;
        RECT 101.530 18.370 101.760 21.150 ;
        RECT 102.320 18.780 102.550 21.370 ;
        RECT 104.000 20.830 104.160 22.420 ;
        RECT 105.860 20.830 106.320 20.835 ;
        RECT 106.650 20.830 107.110 20.835 ;
        RECT 107.440 20.830 107.900 20.835 ;
        RECT 108.230 20.830 108.690 20.835 ;
        RECT 109.020 20.830 109.480 20.835 ;
        RECT 104.000 20.630 109.480 20.830 ;
        RECT 104.000 18.840 104.150 20.630 ;
        RECT 105.860 20.605 106.320 20.630 ;
        RECT 106.650 20.605 107.110 20.630 ;
        RECT 107.440 20.605 107.900 20.630 ;
        RECT 108.230 20.605 108.690 20.630 ;
        RECT 109.020 20.605 109.480 20.630 ;
        RECT 104.000 18.800 105.500 18.840 ;
        RECT 116.200 18.800 116.600 18.890 ;
        RECT 102.320 18.540 103.100 18.780 ;
        RECT 102.320 18.370 102.550 18.540 ;
        RECT 102.910 17.670 103.100 18.540 ;
        RECT 104.000 18.570 107.355 18.800 ;
        RECT 114.405 18.570 116.600 18.800 ;
        RECT 104.000 18.490 105.500 18.570 ;
        RECT 98.480 17.660 103.100 17.670 ;
        RECT 98.480 17.490 103.090 17.660 ;
        RECT 99.910 10.290 100.140 16.090 ;
        RECT 101.550 15.840 101.850 17.490 ;
        RECT 103.400 16.530 103.900 16.540 ;
        RECT 103.400 16.300 109.310 16.530 ;
        RECT 103.400 16.290 103.900 16.300 ;
        RECT 99.900 10.090 100.140 10.290 ;
        RECT 101.570 10.090 101.800 15.840 ;
        RECT 99.900 9.940 100.100 10.090 ;
        RECT 99.400 9.890 102.350 9.940 ;
        RECT 103.400 9.890 103.600 16.290 ;
        RECT 116.200 13.440 116.600 18.570 ;
        RECT 116.200 12.640 149.650 13.440 ;
        RECT 96.170 9.710 96.760 9.725 ;
        RECT 99.400 9.710 103.600 9.890 ;
        RECT 96.110 9.690 103.600 9.710 ;
        RECT 96.110 9.400 99.910 9.690 ;
        RECT 96.110 9.390 98.180 9.400 ;
        RECT 99.400 9.390 99.860 9.400 ;
        RECT 96.170 7.620 96.760 9.390 ;
      LAYER via ;
        RECT 149.320 12.885 149.580 13.145 ;
      LAYER met2 ;
        RECT 149.250 12.640 149.650 13.440 ;
      LAYER via2 ;
        RECT 149.310 12.875 149.590 13.155 ;
      LAYER met3 ;
        RECT 117.850 13.890 149.710 44.290 ;
        RECT 149.250 12.640 149.650 13.890 ;
      LAYER via3 ;
        RECT 149.290 43.730 149.610 44.050 ;
        RECT 149.290 43.330 149.610 43.650 ;
        RECT 149.290 42.930 149.610 43.250 ;
        RECT 149.290 42.530 149.610 42.850 ;
        RECT 149.290 42.130 149.610 42.450 ;
        RECT 149.290 41.730 149.610 42.050 ;
        RECT 149.290 41.330 149.610 41.650 ;
        RECT 149.290 40.930 149.610 41.250 ;
        RECT 149.290 40.530 149.610 40.850 ;
        RECT 149.290 40.130 149.610 40.450 ;
        RECT 149.290 39.730 149.610 40.050 ;
        RECT 149.290 39.330 149.610 39.650 ;
        RECT 149.290 38.930 149.610 39.250 ;
        RECT 149.290 38.530 149.610 38.850 ;
        RECT 149.290 38.130 149.610 38.450 ;
        RECT 149.290 37.730 149.610 38.050 ;
        RECT 149.290 37.330 149.610 37.650 ;
        RECT 149.290 36.930 149.610 37.250 ;
        RECT 149.290 36.530 149.610 36.850 ;
        RECT 149.290 36.130 149.610 36.450 ;
        RECT 149.290 35.730 149.610 36.050 ;
        RECT 149.290 35.330 149.610 35.650 ;
        RECT 149.290 34.930 149.610 35.250 ;
        RECT 149.290 34.530 149.610 34.850 ;
        RECT 149.290 34.130 149.610 34.450 ;
        RECT 149.290 33.730 149.610 34.050 ;
        RECT 149.290 33.330 149.610 33.650 ;
        RECT 149.290 32.930 149.610 33.250 ;
        RECT 149.290 32.530 149.610 32.850 ;
        RECT 149.290 32.130 149.610 32.450 ;
        RECT 149.290 31.730 149.610 32.050 ;
        RECT 149.290 31.330 149.610 31.650 ;
        RECT 149.290 30.930 149.610 31.250 ;
        RECT 149.290 30.530 149.610 30.850 ;
        RECT 149.290 30.130 149.610 30.450 ;
        RECT 149.290 29.730 149.610 30.050 ;
        RECT 149.290 29.330 149.610 29.650 ;
        RECT 149.290 28.930 149.610 29.250 ;
        RECT 149.290 28.530 149.610 28.850 ;
        RECT 149.290 28.130 149.610 28.450 ;
        RECT 149.290 27.730 149.610 28.050 ;
        RECT 149.290 27.330 149.610 27.650 ;
        RECT 149.290 26.930 149.610 27.250 ;
        RECT 149.290 26.530 149.610 26.850 ;
        RECT 149.290 26.130 149.610 26.450 ;
        RECT 149.290 25.730 149.610 26.050 ;
        RECT 149.290 25.330 149.610 25.650 ;
        RECT 149.290 24.930 149.610 25.250 ;
        RECT 149.290 24.530 149.610 24.850 ;
        RECT 149.290 24.130 149.610 24.450 ;
        RECT 149.290 23.730 149.610 24.050 ;
        RECT 149.290 23.330 149.610 23.650 ;
        RECT 149.290 22.930 149.610 23.250 ;
        RECT 149.290 22.530 149.610 22.850 ;
        RECT 149.290 22.130 149.610 22.450 ;
        RECT 149.290 21.730 149.610 22.050 ;
        RECT 149.290 21.330 149.610 21.650 ;
        RECT 149.290 20.930 149.610 21.250 ;
        RECT 149.290 20.530 149.610 20.850 ;
        RECT 149.290 20.130 149.610 20.450 ;
        RECT 149.290 19.730 149.610 20.050 ;
        RECT 149.290 19.330 149.610 19.650 ;
        RECT 149.290 18.930 149.610 19.250 ;
        RECT 149.290 18.530 149.610 18.850 ;
        RECT 149.290 18.130 149.610 18.450 ;
        RECT 149.290 17.730 149.610 18.050 ;
        RECT 149.290 17.330 149.610 17.650 ;
        RECT 149.290 16.930 149.610 17.250 ;
        RECT 149.290 16.530 149.610 16.850 ;
        RECT 149.290 16.130 149.610 16.450 ;
        RECT 149.290 15.730 149.610 16.050 ;
        RECT 149.290 15.330 149.610 15.650 ;
        RECT 149.290 14.930 149.610 15.250 ;
        RECT 149.290 14.530 149.610 14.850 ;
        RECT 149.290 14.130 149.610 14.450 ;
      LAYER met4 ;
        RECT 149.210 13.950 149.690 44.230 ;
  END
END tt_um_Maj_opamp
END LIBRARY

